module grammer

pub const reserved_symbols = {
	'import':     ['prayog']
	'as':         ['naam']
	'false':      ['bethik']
	'true':       ['thik']
	'function':   ['karya']
	'if':         ['yedi']
	'else':       ['natra']
	'loop':       ['ghum', 'for']
	'break':      ['todh']
	'continue':   ['xod']
	'return':     ['pathau']
	'nil':        ['khali', 'null', 'sunna']
	'v':          []
	'endv':       []
	'del':        ['hatau']
	'__module__': []
	// predefined functions
	'assert':     ['pariksan']
	'panic':      ['truti']
	'print':      ['dekhau']
	'println':    ['dekhauln']
	'input':      ['sodha']
	'len':        ['ginti']
	'typeof':     ['prakar']
	'int':        ['aanka']
	'table':      []
	'float':      []
	'string':     ['sabda']
	'chr':        []
	'rand_str':   []
	'rand_int':   []
	'server':   []
	// 'not':      ['hoina']
	// 'or':       ['ya']
	// 'and':      ['ra']
}
