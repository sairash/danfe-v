module parser

import lexer

pub struct Parse {
	mut:
		lex *lexer.Lex
}

