module grammer

pub const reserved_symbols = [
	'false',
	'true',
	'function',
	'if',
	'else',
	'loop',
	'break',
	'print',
	'input',
	'nil',
	'not',
	'or',
]
