module grammer

pub const reserved_symbols = {
	'import':   ['ayat', 'prayog', 'include']
	'as':       ['naam']
	'false':    ['bethik']
	'true':     ['thik']
	'function': ['karya', 'func']
	'if':       ['yedi']
	'else':     ['natra', 'fi']
	'loop':     ['ghum', 'for', 'while', 'until']
	'break':    ['todh']
	'continue': ['xod']
	'return':   ['pathau']
	'print':    ['dekhau']
	'println':  ['dekhauln']
	'input':    ['sodha']
	'nil':      ['khali', 'null', 'sunna']
	// 'not':      ['hoina']
	// 'or':       ['ya']
	// 'and':      ['ra']
}
