module grammer

pub const reserved_symbols = {
	'import':     ['ayat', 'prayog', 'include']
	'as':         ['naam']
	'false':      ['bethik']
	'true':       ['thik']
	'function':   ['karya', 'func']
	'if':         ['yedi']
	'else':       ['natra']
	'loop':       ['ghum', 'for', 'while', 'until']
	'break':      ['todh']
	'continue':   ['xod']
	'return':     ['pathau']
	'nil':        ['khali', 'null', 'sunna']
	'v':          []
	'endv':       []
	'del':        ['hatau']
	'__module__': []
	// predefined functions
	'print':      ['dekhau']
	'println':    ['dekhauln']
	'input':      ['sodha']
	'len':        ['ginti']
	'typeof':     ['prakar']
	'push':       ['hala']
	'pop':        ['nikala']
	// 'not':      ['hoina']
	// 'or':       ['ya']
	// 'and':      ['ra']
}
